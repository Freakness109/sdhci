// Copyright 2025 ETH Zurich and University of Bologna.
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51

// Authors:
// - Micha Wehrli <miwehrli@student.ethz.ch>
// - Axel Vanoni <axvanoni@student.ethz.ch>

module tb_acmd12 #(
    parameter time         ClkPeriod     = 50ns,
    parameter int unsigned RstCycles     = 1
  )();

  int ClkEnPeriod;

  sdhci_fixture #(
    .ClkPeriod(ClkPeriod),
    .RstCycles(RstCycles)
  ) fixture ();

  // < 0 cmd12 gets delayed due to our command
  // = 0 both requests arrive at the same time, cmd12 goes first
  // > 0 our command gets delayed by cmd12
  int CyclesThatDriverCommandArrivesBeforeCMD12;
  int IsFirstResponseValid;

  logic AutoCMD12First;
  logic [15:0] normal_status;
  logic [15:0] error_status;
  logic [15:0] cmd12_error_status;
  logic cmd_en;
  logic dat_en;

  initial begin
    $timeformat(-9, 0, "ns", 12);
    $dumpfile("tb_acmd12.vcd");
    $dumpvars(0);

    if (!$value$plusargs("CyclesThatDriverCommandArrivesBeforeCMD12=%d", CyclesThatDriverCommandArrivesBeforeCMD12)) begin
      CyclesThatDriverCommandArrivesBeforeCMD12 = 0;
    end
    if (!$value$plusargs("IsFirstResponseValid=%d", IsFirstResponseValid)) begin
      IsFirstResponseValid = 0;
    end
    if (!$value$plusargs("ClkEnPeriod=%d", ClkEnPeriod)) begin
      ClkEnPeriod = 4;
    end

    AutoCMD12First = CyclesThatDriverCommandArrivesBeforeCMD12 <= 0;

    $display("Testing auto cmd12 with CyclesThatDriverCommandArrivesBeforeCMD12=%d, IsFirstResponseValid=%d, ClkEnPeriod=%d", CyclesThatDriverCommandArrivesBeforeCMD12, IsFirstResponseValid, ClkEnPeriod);

    fixture.vip.wait_for_reset();

    fixture.vip.set_interrupt_status_enable(
      .normal_interrupt_status_enable('hFFFF),
      .error_interrupt_status_enable('hFFFF),
      .finish_transaction(1'b0)
    );

    fixture.vip.set_frequency_select(
      .divider(8'(ClkEnPeriod >> 1)),
      .finish_transaction(1'b0)
    );

    fixture.vip.set_clock_enable(.enable(1'b1), .finish_transaction(1'b0));

    fixture.vip.set_transfer_mode(
      .is_multi_block(1'b0),
      .is_read(1'b0),
      .auto_cmd12_enable(1'b1),
      .block_count_enable(1'b1),
      .dma_enable(1'b0),
      .finish_transaction(1'b0)
    );

    fixture.vip.set_block_size_count(
      .block_size(12'd64),
      .block_count(16'd1),
      .finish_transaction(1'b0)
    );

    fixture.vip.launch_command(
      .command_index(6'd0),
      .command_type (2'b00), // normal command
      .data_present (1'b1),
      // no response -> no checking
      .index_check_enable(1'b0),
      .crc_check_enable(1'b0),
      .response_type(2'b00), // no response
      .finish_transaction(1'b1)
    );

    repeat(10) fixture.vip.wait_for_sdclk();
    repeat (64 / 4) begin
      fixture.vip.write_buffer_data('hDEAD_BEEF);
      fixture.vip.wait_for_sdclk();
    end


    // These values are slightly random because of the offset between command start and sd clk period
    case (ClkEnPeriod)
      1: repeat(539 - CyclesThatDriverCommandArrivesBeforeCMD12) fixture.vip.wait_for_clk();
      2: repeat(1077 - CyclesThatDriverCommandArrivesBeforeCMD12) fixture.vip.wait_for_clk();
      4: repeat(2155 - CyclesThatDriverCommandArrivesBeforeCMD12) fixture.vip.wait_for_clk();
      default: $fatal("ClkEnPeriod not supported");
    endcase

    fixture.vip.launch_command(
      .command_index(6'd0),
      .command_type (2'b00), // normal command
      .data_present (1'b0),
      .index_check_enable(1'b1),
      .crc_check_enable(1'b1),
      .response_type(2'b10) // 48bit no busy
    );

    fixture.vip.wait_for_sdclk();
    repeat(80) fixture.vip.wait_for_sdclk();

    if (IsFirstResponseValid) begin
      // valid response, next command should run
      if (AutoCMD12First)
        fixture.vip.send_response_48(12, 'h7A);
      else
        fixture.vip.send_response_48(0, '0);
    end else
      // invalid response, next command should not run
      fixture.vip.send_response_48('1, '1);

    if (IsFirstResponseValid) begin
      repeat(80) fixture.vip.wait_for_sdclk();

      // Valid response for the second command
      if (AutoCMD12First) begin
        fixture.vip.send_response_48(0, '0);
      end else begin
        fixture.vip.send_response_48(12, 'h7A);
      end
    end else begin
      repeat (80*ClkEnPeriod) begin
        // TODO: make a wait for command
        fixture.vip.wait_for_clk();
        fixture.vip.test_delay();
        fixture.vip.is_cmd_held(cmd_en);
        if (cmd_en) $fatal("Second command should not have been sent");
      end
    end

    repeat(10) fixture.vip.wait_for_sdclk();

    fixture.vip.get_interrupt_status(
      .normal_interrupt_status(normal_status),
      .error_interrupt_status(error_status)
    );
    error_status[15:4] = '0; // Only care about cmd errors

    fixture.vip.get_acmd_error_status(cmd12_error_status);

    // leave some time so we get a cleaner waveform
    repeat(10) fixture.vip.wait_for_clk();

    if (IsFirstResponseValid) begin
      if (|(error_status)) begin
        $error("Got an error when we shouldnt have 0x%h", error_status);
        $fatal();
      end
      if (|(cmd12_error_status)) begin
        $error("Got a cmd12 error when we shouldnt have 0x%h", cmd12_error_status);
        $fatal();
      end
    end else begin
      if (AutoCMD12First) begin
        if (|(error_status)) begin
          $error("Got an error when we shouldnt have 0x%h", error_status);
          $fatal();
        end
        if (cmd12_error_status != /* command not issues by acmd12 error + crc error + index error */ 'b1001_0100) begin
          $error("Got a cmd12 error when we shouldnt have 0x%h", cmd12_error_status);
          $fatal();
        end
      end else begin
        if (error_status != /* crc error + index error */ 'b1010) begin
          $error("Got an error when we shouldnt have 0x%h", error_status);
          $fatal();
        end
        if (cmd12_error_status != /* command not executed */ 'b1) begin
          $error("Got a cmd12 error when we shouldnt have 0x%h", cmd12_error_status);
          $fatal();
        end
      end
    end

    $dumpflush;
    $finish();
  end

endmodule
