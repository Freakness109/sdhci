module sd_bus_dat_driver (
  input   logic dat0_i,
  input   logic dat1_i,
  input   logic dat2_i,
  input   logic dat3_i,

  input   logic dat_highz_i,
  input   logic dat0_pull_up_i
);
  
endmodule