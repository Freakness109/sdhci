module sd_bus_cmd_receiver (
  output  logic cmd_o
);
  //hook up to cmd line
  assign cmd_o = 0'b0;
endmodule